library verilog;
use verilog.vl_types.all;
entity barrelShifter_tb is
end barrelShifter_tb;
