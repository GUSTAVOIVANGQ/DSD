library verilog;
use verilog.vl_types.all;
entity FDD_FPGA_tb is
end FDD_FPGA_tb;
