library verilog;
use verilog.vl_types.all;
entity FFJK_tb is
end FFJK_tb;
