library verilog;
use verilog.vl_types.all;
entity tb_jk_bcd is
end tb_jk_bcd;
